`ifndef MY_CASE0__SV
`define MY_CASE0__SV

class long_seq extends uvm_sequence#(my_transaction);
    // rand bit[47:0] dmac; //name collision!!!
    rand bit[47:0] ldmac; 
    `uvm_object_utils(long_seq)
    function  new(string name= "long_seq");
        super.new(name);
    endfunction 
    
    virtual task body();
        my_transaction tr;
        `uvm_do_with(tr, { tr.crc_err == 0;
                           tr.pload.size() == 1500;
                           tr.dmac == ldmac;})
        tr.print();
    endtask
endclass

class case0_sequence extends uvm_sequence #(my_transaction);

    function  new(string name= "case0_sequence");
        super.new(name);
        set_automatic_phase_objection(1);
    endfunction
   
    virtual task body();
        long_seq lseq;
        repeat (10) begin
            `uvm_do_with(lseq, {lseq.ldmac == 48'hFFFF;})
        end
        #100;
   endtask

   `uvm_object_utils(case0_sequence)
endclass

class my_case0 extends base_test;

    function new(string name = "my_case0", uvm_component parent = null);
        super.new(name,parent);
    endfunction 
    extern virtual function void build_phase(uvm_phase phase); 

    `uvm_component_utils(my_case0)
endclass


function void my_case0::build_phase(uvm_phase phase);
    super.build_phase(phase);

    uvm_config_db#(uvm_object_wrapper)::set(
        this, 
        "env.i_agt.sqr.main_phase", 
        "default_sequence", 
        case0_sequence::type_id::get()
    );
endfunction

`endif
