`ifndef MY_CASE0__SV
`define MY_CASE0__SV

class sequence0 extends uvm_sequence #(my_transaction);
    my_transaction m_trans;

    function  new(string name= "sequence0");
        super.new(name);
        set_automatic_phase_objection(1);
    endfunction

    virtual task body();
        repeat (2) begin
            `uvm_do(m_trans)
            `uvm_info("sequence0", "send one transaction", UVM_MEDIUM)
        end

        // 鎖死 1st
        lock();
        `uvm_info("sequence0", "locked the sequencer ", UVM_MEDIUM)
        repeat (5) begin
            `uvm_do(m_trans)
            `uvm_info("sequence0", "send one transaction", UVM_MEDIUM)
        end
        `uvm_info("sequence0", "unlocked the sequencer ", UVM_MEDIUM)
        unlock();

        repeat (2) begin
            `uvm_do(m_trans)
            `uvm_info("sequence0", "send one transaction", UVM_MEDIUM)
        end
        #100;
    endtask

    `uvm_object_utils(sequence0)
endclass

// second seq
class sequence1 extends uvm_sequence #(my_transaction);
    my_transaction m_trans;

    function  new(string name= "sequence1");
        super.new(name);
        set_automatic_phase_objection(1);
    endfunction

    virtual task body();
        repeat (3) begin
            `uvm_do_with(m_trans, {m_trans.pload.size < 500;})
            `uvm_info("sequence1", "send one transaction", UVM_MEDIUM)
        end

        // 鎖死 2nd
        lock();
        `uvm_info("sequence1", "locked the sequencer ", UVM_MEDIUM)
        repeat (4) begin
            `uvm_do_with(m_trans, {m_trans.pload.size < 500;})
            `uvm_info("sequence1", "send one transaction", UVM_MEDIUM)
        end
        `uvm_info("sequence1", "unlocked the sequencer ", UVM_MEDIUM)
        unlock();

        repeat (3) begin
            `uvm_do_with(m_trans, {m_trans.pload.size < 500;})
            `uvm_info("sequence1", "send one transaction", UVM_MEDIUM)
        end
        #100;
    endtask

    `uvm_object_utils(sequence1)
endclass

class my_case0 extends base_test;

    function new(string name = "my_case0", uvm_component parent = null);
        super.new(name,parent);
    endfunction 
    extern virtual task main_phase(uvm_phase phase);

    `uvm_component_utils(my_case0)
endclass


task my_case0::main_phase(uvm_phase phase);
    sequence0 seq0;
    sequence1 seq1;

    seq0 = new("seq0");
    seq0.starting_phase = phase;
    seq1 = new("seq1");
    seq1.starting_phase = phase;
    fork
        seq0.start(env.i_agt.sqr);
        seq1.start(env.i_agt.sqr);
    join

endtask

`endif
