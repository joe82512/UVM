`ifndef A_BLOCK_TRANSPORT__SV
`define A_BLOCK_TRANSPORT__SV

class A extends uvm_component;
    `uvm_component_utils(A)

    uvm_blocking_transport_port#(my_transaction, my_transaction) A_transport;
    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction

    extern function void build_phase(uvm_phase phase);
    extern virtual  task main_phase(uvm_phase phase);
endclass

function void A::build_phase(uvm_phase phase);
    super.build_phase(phase);
    A_transport = new("A_transport", this);
endfunction

task A::main_phase(uvm_phase phase);
    my_transaction tr;
    my_transaction rsp;
    repeat(10) begin
        #10;
        tr = new("tr");
        assert(tr.randomize());
        A_transport.transport(tr, rsp);
        `uvm_info("A", "received rsp", UVM_MEDIUM)
        rsp.print();
    end
endtask

`endif
